typedef uvm_sequencer #(alu_tx) alu_sequencer;


